-------------------------------------------------------------------------------
--
-- Title       : top_tb
-- Design      : range_finder
-- Author      : Michal
-- Company     : AGH
--
-------------------------------------------------------------------------------
--
-- File        : C:\My_Designs\project_PSC\range_finder\src\top_tb.vhd
-- Generated   : Fri Jan  3 20:03:51 1992
-- From        : interface description file
-- By          : Itf2Vhdl ver. 1.22
--
-------------------------------------------------------------------------------
--
-- Description : 
--
-------------------------------------------------------------------------------

--{{ Section below this comment is automatically maintained
--   and may be overwritten
--{entity {top_tb} architecture {top_tb}}



entity top_tb is
end top_tb;

--}} End of automatically maintained section

architecture top_tb of top_tb is
begin

	 -- enter your statements here --

end top_tb;
